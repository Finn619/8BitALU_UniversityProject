library verilog;
use verilog.vl_types.all;
entity Multi21_vlg_vec_tst is
end Multi21_vlg_vec_tst;
