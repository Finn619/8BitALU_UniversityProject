library verilog;
use verilog.vl_types.all;
entity ShiftingUnit_vlg_vec_tst is
end ShiftingUnit_vlg_vec_tst;
