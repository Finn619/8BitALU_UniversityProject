library verilog;
use verilog.vl_types.all;
entity CLAAdder_vlg_vec_tst is
end CLAAdder_vlg_vec_tst;
