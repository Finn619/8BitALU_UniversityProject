library verilog;
use verilog.vl_types.all;
entity LogicUnit_vlg_vec_tst is
end LogicUnit_vlg_vec_tst;
