library verilog;
use verilog.vl_types.all;
entity Multi21 is
    port(
        Y               : out    vl_logic;
        pin_name1       : in     vl_logic;
        I1              : in     vl_logic;
        I0              : in     vl_logic
    );
end Multi21;
